        ?  &�      �  h      ,                  �    NV��B���J� m&�    l .  |  ?(/0 /<  Zva�    POB����   ���dD".�� ЀЁЀ |  ?h���   ��� fP ЀЁЀ |  ?i���   ��� f2R���J���g$".�� ЀЁЀ |  ?j��//<  Z�a�    PON^NuR���` �~NV  /.. J�    g@ r��   ��   �g � ���� ���f/<  �/<  Z�/<  Z�a�    �� J�    gD r��   ���    g0 r��   ���    g/<  �/<  [/<  Z�a�    �� J�    g0 r��   ��    e/<  �/<  [?/<  [a�    �� J�    g4 r��   � |    J� f/<  �/<  [r/<  [Pa�    �� J�    gB r��   � |     p  ���   �J� f/<  �/<  [�/<  [�a�    �� J�    gP r��   � |     p  ���   � p  ��   J� f/<  �/<  \/<  [�a�    ��  r��   � |     p  ���   � p  ��    0 .N^NuNV  //*n ~ `:p /  L|   J�g <  \/`
     <  \1/ /<  \(a�    �� R��� m�/<  \4a�    XO.*_N^NuNV�� n /( (a�����XO-@�� 9    �   �g/<  \6a�    XO n  �    n��( I�r� n !A  n !A `"n  I"i @#h  HB�/<    n r��( Jf n�� ( Ё`       n ( JI�/  n  ( (��   / /<   (/. a�    �� N^NuNV��/////*n (n ~ | &L�� � K-|  \F�� , �   @f  � , �   �g  ���   f
+ ( g  �r)�+ fJ+ f/- (/<  \Ga�    `  �     l �/( /- d/- (/<  \�a�    ��  l �//<  \�a�    POp + / p + / �� �   �/ /<  \�a�    �� �� g/+ /<  \�a�    PO/<  ]a�    XO/<  ]	a�    XO - �� `/ /a�����PO�  �� G  qf  ���   f/<  ]$a�    XOR�`  �    �� � [ f/<  ]:a�    XO~`  �  /<  ]Wa�    XOp + / �� �   �/ /<  ]{a�    �� /<  ]�a�    XO`T    �� �   �@ b � p�  �N�    �  X  p  @  p  p  �  p  p  p  �  �J�g4 , �   @f(p + / p + / �� �   �/ a������� J�f �   g B| ` B  ~ l ��   g�-|  ]��� , �   @f ���� g ��/<  ]�/.��/<  ]�a�    �� /+  - (� ���/ /<  ]�a�    �� ` �F    R�` �<  p + @ (b  �g(J@g �$@ g �@ g �@ g �~` �
    �  - M  J g �   g~` ��      - MI��  @ M0- NH��  ;@ N l ������p��� �����R�` ��@ )g�@ *g ��@ Gg�@ Hg�` �z  ~` ��   �    ;@ $g �    ,.&_(_*_N^NuNV  ///*n /- (a����XO(@&L�� � K 9    �  �g"/+ p + / p / /<  ]�a�    ��  9    �  �gp / Hk a�����PO+k  </<   B�p / Hk /a�    �� &_(_*_N^NuNV  //*n /- (/<  ^6a�    PO/a�    XO(m @ m 0 (  �   gN�   !|  >J� :g
 l : �    J, CfN|  AB� m 0( (I�/ //<    Hl ,a�    �� `"J, Cg�J� :f|  >`     l : �    (_*_N^NuNV  //*n  m @( AI�/ /- (/<  ^^a�    �� (m @ m 0 (  �   gN�   !|  >J� :g
 l : �    J, CfN|  AB� m 0( (I�/ //<    Hl ,a�    �� `"J, Cg�J� :f|  >`     l : �    (_*_N^NuNV  //*n /- (/<  ^�a�    PO/a�    XO(m @ m 0 (  �   gR�   !|  >J� :g
 l : �    J, CfR|  AB� m 0( (I�/ //<    Hl ,a�    �� `&    J, Cg�J� :f|  >`     l : �    (_*_N^NuNV  /*n B� m 0( (I�/ //<    /- (a����4XO�  4/ a�    �� *_N^NuNV��////
//*n (m @/- (a�����XO&@a�    J�g zHn��a�    XOB� :B, >rA C�� 0e  � 9    �   g, AI�/ /- (/<  ^�a�    �� Hl a�    XOJ, >gB, >/<   a�    XO, AH�@ n �g �@ n �g  �J@g@ gU@gL` HB� d|  A/<  
�/a�    POB, CJ, >gB, >/<   a�    XOHn��a�    ` z    B, BB- IHl /9  ?//<  	�a�    �� �����/a�    XO. g�Hl a�    XOJ, >gB, >/<   a�    XOU�f �r 9    �   g �R- KI�/ /<  ^�a�    PO` �8    | 
 A/a�    XO �   ;|  $ 9    �   g/- (/<  ^�a�    PO �   g�����/a�    XO/a�    XO` ��    /- (/<  _a�    PO/<   a�    XO/a�    XO �   B, A` �/<   a�    XO|  A �   |  I �   f �x` �d/a�    XOJ�g ��//<  
ba�    ` �P       9    �   g �/<  _"a�    XO` �       9    �   g �/<  _?a�    XO` �       9    �   g �/<  _Za�    XO` �      ����� 9    �   g/<  _oa�    XO|  L/<  
�/a�    POHl /- <//<  >a�    �� ` 8   9    �   g/<  _�a�    XO0- N@ J@g@0- NH��  ;@ N k � �   B� \ 9    �   g 
�/<  _�a�    XO` 
�   9    �   g 
�/- (/<  _�a�    PO` 
�  J+Fm2 +BF���    �     8f  - �� H�+FI� |    Ѱ ����� 9    �   g/<  _�a�    XO, B  J g, B  J f"/<  `/<  `a�    PO/<   a�    XOJ- Lg 
J� `g6 k �+h   k �*�+l ` ,B� `/<  `$a�    XO/<   a�    XO-  Lf`)m , ` K�� �+H , k �!m   k �!m `  k � � k �!m 8  �   |  A+|     8` �(    �     8f ��` ��-  LfP , dR� d��  ?l8/a�    XO|  A �   B�/<   2//<  
ba�    �� ` 	    ;|  $`;|  $ �   J� `g  �+l ` ,B� `�     8g/<  `Aa�    XO k �+h  8 k �*��� �U f  � , dR� d��  ?l/a�    XO|  A k �+h  ` �R;|  $ �   �� �@ M k �+h  ` k �+h  | 
 A/a�    XOJm $g* �    9    �   g0- $H�/ /<  `_a�    PO/a�    XO` //a����POJ�g ��|  A k �+h   k �+h  ` �   ` ��   9    �   g/<  `sa�    XOS�R��   �. ��l
| ` �    S�S�R� f �0- N@ J@g vR�Z��R��U�B� \p2�.��b  �p .��@ �b  �J.��g  �p�.��cp .���)@ \p .��@ �cp `  ~      p}�.��d <   �`  f      pd�.��d <   �`  N      p^�.��d <  �`6pK�.��d <   �`&p?�.��d <  �`p2�.��d <   �` <  ��� \J+FmVJ.��gP/9  ?/9  ?p .��/ a�    XO// a�    �� -A��-@��//.��a�    PO+FI� |    !�  k � �   0- NH��  ;@ N 9    �   g 0/, \/<  `�a�    PO`     /<  `�a�    XO V�/ Hj��a����VPO�ǜ�` �p @ �J@g, 9    �   g �p / /<  `�a�    PO` �    p / /<  `�a�    PO/<   a�    XO` �   �   g ��` �,| J- If  �J+FmJ +B��    �     8f,+FI� |    R� +FI� |    R� `  r@`,    �     8g� - (��   �   �"�   f�r Ё�h�R� �   g� h�R�`  x   k � �0   �    f`B� \Hvh�/a�    PO. ܇�   fB0- NH��  ;@ N`2      0- N@ J@g � h�R�0- NH�� ;@ NB� \�����J�f� h�R������|  IHl /9  ? //<  �a�    �� /Hn��/a�    �� Hl a�    XOJ, >gB, >/<   a�    XO �   g�����/<   a�    XO|  A` ��  |  IJ, Bg$/<  a/<  aa�    PO/<   a�    XO`, BI��  @ B)m  H)m , DHl /9  ? //<  �a�    �� / m 8N�XO` ��    /<  a2/<  a!a�    PO/<   a�    XO|  I 9    �   g/, D/, H/<  a@a�    �� Hl /9  ? //<  �a�    ��  �   g& m 0( %�   �/ a�    XOJ�f
�     8f./<    �   / /, H/, D/a�    �� ` ��      �     8g�/<   `�      , B  J f, BI�� @ B`&    /<  au/<  ada�    PO/<   a�    XO|  I m @ - �� H�� `Hl /9  ? //<  �a�    �� /a�    XO@ L  �g|  AHl a�    XOJ, >gB, >/<   a�    XOJ- Lg �z 9    �   g �j- LI�/ /<  a�a�    PO` �P    /<   a�    XO�����- II�/ , AI�/ /<  a�a�    �� , BI�/ /<  a�a�    PO/<   a�    XO` �    @ g ��@ g ��]@f�` ��@ An:g@ g ��@ 	g �r@ @f �x, B  J g ��, BI�� @ B` ��@ Bg �@ Cg �R@ Fg �R@ Gf �8 �   g �   Hl /9  ? //<  �a�    �� Hn��/a�    PO, Hl a�    XOJ, >gB, >/<   a�    XO|  A$N���� Jp�- IfS�R�|  I S�J�g ��p @ b �D p�  (N�  �  p  H  p  �  `  `    �R�`�Hl a�    XOB, > |  //- (/<  a�a�    �� /- /- d/<  b	a�    �� J+Fm +BF���    /a�    XO| 
 AB� `/a�    XOJ�g/- (/<  b(a�    PO/a�    XO �   f2 |  �   g$�   g�   g �   B, A` �       �   ;|  $/a�    XO,.$_&_(_*_N^NuNV  /. a�    XON^NuNV  ///*n (n /- (a����JXO&@ �   �����Bm $ - (r��   � |    +p  0k  H - (���   �@ K+|  
� 4B- J+|  .� < +@ D . �   b  � p�  �N�     H  X  p  0  �  �//+ �a�    PO&_(_*_N^NuB� <+|  F 4`�  l  J+|  � <+|     8`�+|     8`�      B� D+|  FP <+|     8`�  l  JB� D+|  FP <+|     8` �|  +|     8` �n    +|     8` �^    /<  bPa�    XO` �HNV��//*n �     f/<   �a�    XO(@`X       9    �   gr��    /9    a�    XO`�  r��    J�    f/<   �a�    XO#�    (y    (�   J�  g
 �   `  ���������� � �  B, MBl N)n  (Bl $n ' J . r��   � |    )p  0 . ���   �@ Km  H)n  <)n  4)n  8B� D�     f. '�   �/ /, ,/. a�    �� //- �a�    PO/a�    XO �   f  tJ� g&�     g , �� `/ /. /, ,a�    �� �     f< , �� `@  9    �   g"/<  bla�    XO- I�/ Hm a����(PO�     f  �B� B-  �   f  �J� `f  �J� `f  |/<   Hm /, ,a�    �� /<   Hn�� l ,Hh a�    �� R�  9    �   g(/.��/- /, (/<  b�a�    �� `
      R-  .���-@��f��     f/a�    XO`$   9    �   g/9    a�    XOB�    /a�    XO(_*_N^NuNV��/////..  r��   � |    *p  f x r��   � |    z�!� -|   `��a�    * -|    �� n��R�  ( S�f n��!E   y    B� n��J�fN y     �   -|    �� n��S� f n��/(  a�    XOB�/<   /<   $a�    �� *@`  �  -|  ��� n��*P � n��R�  n��S�  n��R�  n��R�  n��r@Ө "n�� I (  �� n (  n��!@   y     �   -|    �� n��S� f n��/(  a�    XO r��   ��"<    Ҁ/a�    XO/<   $/a�    PO r��   � |    !� `@    ����f6 r��   ��"<    Ҁ/a�    XO r��   � |    *p  ���   �(u  f j ���   �z�+� -|   ���a�    * -|    �� n��R�  ( S�f n��!E   y    B� n��J�fP y     �   -|    �� n��S� f n��/(  a�    XOB�/<   /<   �a�    �� (@`  �    -|  ��� n��(P � n��R�  n��S�  n��R�  n��R�  n���    "n�� I (  �� n (  n��!@   y     �   -|    �� n��S� f n��/(  a�    XO ���   ��"Ҁ/a�    XO/<   �/a�    PO ���   �+� R�  `2    ����f( ���   ��"Ҁ/a�    XO ���   �(u  ��   &t  f x ��   z�)� -|   ���a�    * -|    �� n��R�  ( S�f n��!E   y    B� n��J�fN y     �   -|    �� n��S� f n��/(  a�    XOB�/<   /<  Ha�    �� &@`  �  -|  ��� n��&P � n��R�  n��S�  n��R�  n��R�  n���    "n�� I (  �� n (  n��!@   y     �   -|    �� n��S� f n��/(  a�    XO ��   �"Ҁ/a�    XO/<  H/a�    PO ��   )� R�   L�� $'H � L�� �'H �`.����f( ��   �"Ҁ/a�    XO ��   &t  R�J�f � ���'@ | �F *.&_(_*_N^NuNV��/////.. �͙̗� r��   � |    *p  g � ���   �(u  g � ��   &t  g xS�f r + �   g
z�˫ ` \ ��   B� S�  /a�    XO-@��J�    g, / a�    XOJ�f/<  �/<  d/<  c�a�    ��  n��P c/<   /a�    PO`  �       n��0�  ��� |    ��-H��-|  ���J�    g& n��Jh g/<  �/<  d+/<  da�    �� a�    * -|    �� n��R�  ( S�f n��!E   y    B� n��&� n�� � n��S�  n��0�  ��r� n����  n��R�  y     �   -|    �� n��S� f n��/(  a�    XO g dJ�  f \ ���   �B� S�  /a�    XO-@��J�    g, / a�    XOJ�f/<  �/<  d�/<  d_a�    ��  n��P c/<   /a�    PO`  �       n��0�  ��� |    ��-H��-|  ���J�    g& n��Jh g/<  �/<  d�/<  d�a�    �� a�    * -|    �� n��R�  ( S�f n��!E   y    B� n��(� n�� � n��S�  n��0�  ��r� n����  n��R�  y     �   -|    �� n��S� f n��/(  a�    XO g dJ�  f \ r��   � |    B� /a�    XO-@��J�    g, / a�    XOJ�f/<  �/<  d�/<  d�a�    ��  n��P c/<   /a�    PO`  �   n��0�  ��� |    ��-H��-|  ���J�    g& n��Jh g/<  �/<  e#/<  ea�    �� a�    * -|    �� n��R�  ( S�f n��!E   y    B� n��*� n�� � n��S�  n��0�  ��r� n����  n��R�  y     �   -|    �� n��S� f n��/(  a�    XO*.&_(_*_N^NuNV  //..  �   g/a�    XO.*_N^Nu/a�����XO*@�   gJ�  C�g&B�/<   /<   �B�/B�/<  F/a�������  �   f</a�  XO�   ��  gr�í  r��   � |    /0 a�    XO r��   ���    fS� fHr�í `@ �� �   f2��  g*B�/<   /<   �B�//<    /<  
�/a����"��  /a����<XOp ` �NV  ////..  �   g/. /a�    PO,.(_*_N^Nu r��   ��    lR r��   � |    *p  g8p�- $f0 ���   �Q�l" ���   �- &I���g ��   Q�mp` ��/a���� XO(@ fp` �t   , �   f � ����� g/a����ZXOp` �H       r��   ���    f , �   f�R� /a�  �XO�   f  �/a�    XOB�/<   /<   �Hl //<    /<  
�/a������  , g/a�����XO ` ��      /<   /<  e4Hl a�    �� J�fJ/<   /<  e=Hl &a�    �� J�g/<   /<  eNHl &a�    �� J�fr�� `       l � �     r��   ���    fJ �� �   f<�� � �   �@ b* p�  +�N�  ,  ,z  ,z  ,z  ,  ,  ,z  ,~�� p ` ��    B�/<   /<   �B�//<    /<  
�/a������  , f ��/a�  0XO, f ����  g�B�/<   /<   �B�//<    /<  
�/a����P��  ` �|NV  /"n J)Fl  z~ �   l  n |    J�| ffGFp�#@BF���     |    B�|  |    B�|  |    B�|  |    !�  ?|  9    r�") � pҀ |    !�| .N^NuR�` ��NV  "n J)Fm)FI� |    B� | �FN^NuNV��///////*n (n &n /<   /<   /<   2Hn��/. /<    /<  
�/a����>��  . g (*,.&_(_*_N^Nu/<   Hn��a�    PO/<    Hn��Hn��a�    �� | �� gJ�fp 0.��,  g
(�`    , gJ�fp 0.��( `    ( g&�0.���  ���� ��  ���   fr`�   fr	`    rL  * =F��E��=D��/<   $/<   /<   2Hn��/. /<    /<  
�/a����D��  . f � L �+@ �   fp`    �   fp	`    p
@ ` ��NV��////.. *n B���|P-F��Hn��Hn��//a����N�� * g*,.*_N^Nu,.��B�/<   /<  �B�//<  /<  
�/a������  J�g  �-|   ������gFB�Hn��//a������� J�f.B�/<   /<  �B�//<  /<  
�/a����@��  J�g4�   ��f <   `�   ��f <   `      p -@��f ��J���g  �/<����/<   /<  �B�//<  /<  
�/a�������  J�gV|M-F��Hn��Hn��//a����,�� J�f2/<����/<   /<  �B�//<  /<  
�/a������  J�gB���J���gJ���fB� B- p ` ��NV  //. a����DXO*@ - �   g2J� f,B�/<   /<   �B�/. /<    /<  
�/a������   - �   fZr��  - �   gr@�� //. a�����POp��� `,B�/<   /<   �B�/. /<    /<  
�/a������  J� fp*_N^Nup `�NV��/// . �   g �/. /. /. /. a�    �� ` �    g v�  Deg �  Dfg  ��  Dgg ��  Sg�  Sg>p` N.. �?�  r�- I���l- I�//. Hm a�    �� `    - �   g< - �   f/. a����nXO n  � - I�r� n !A ` �      /. a����>XO. g�` �    /. a����&XO. f �- I�"- �p
J�jD��D�`    �S� n  �` v   . �   fa�    J�f
p` Z    �   gp` H   n �   f~�� ` .  ~�ϭ ` "       n J�g�p`    . �   fa�    J�f
p` �    ~�� gp` �   n J�g~�� ` �      ~�ϭ ` �       - �   fp` �       n �   �. �   g�   
g�   g
p` r    /<   Hm �/. a�    �� ` P     . �?�  r��   �d . �?�  r�`   <   �. //. Hm �a�    �� /<   �Hm �a�    PO` �       . �   fa�    J�f
p` �     - �   g  � n 0@ b  � p�  4PN�    4�  4�  4�  4�  4�  5   5   5   5   5   5   5   5   5   5   5   4�Hn��Hn��//. a������� . g  X` @  -|   ��~M-G��`�-|   ��~M-G��`�-|   ��~M-G��`�-|   ��~P-G��` ��      p` �   - �   f$ - �   g�   f~�� `
p` �  ~  n 0( H�/ /<   /< ~@B�/. /<    /<  
�/a����Z��  , S�f~�ϭ  ` t      /<   /<   /<   2Hn��/. /<    /<  
�/a������  -@��.��  J gp`  p  n  � .��`  - �   g,B�/<   /<   �B�/. /<    /<  
�/a������   - �    gp`p  n  �~�ϭ `  �      /<   /. Hm &a�    ��  n r!A /. a����XOJ�g n B�  n B� `$     - S� n !@ - I�r� n !A �� � �   �. fp `.    �   fp`    �   fp`    _�fp`p� n !@ p ,.*_N^Nu/. a���ɸXO*@ . �  ���  So �R�  Sg ��  Sg ���  Sg �l�  Sg �B�  S*g ��` �NNV  ///*n .- (J�    g& �   g/<  �/<  ew/<  e_a�    ��  �   gB�/a�    ` ,  /a����XO(@ r��   � |    +p  0 ���   �@ K�����B- MBm N+y  ?$ <+|  
� 4 r��   ���    f4 , �   g(J, �g
 �   `  �����+|  � 8+m  ``  t/a���� XOJ�g;|  $ �   /a�    XO`  ll  HB�, I�/ /, /a�    �� J�fF �    - (�   g
 <    `   <    +@ 8p 9    � �    //, �a�    PO.(_*_N^NuNV   . �   g/. /. a�    PON^Nu/. /<    B�/. B�/<  7Va�    �� `�NV   . �   g/. /. a�    PON^Nu/. /<    /<   /. B�/<  7Va�    �� `�NV�� . �   g$/. a�    XON^Nu/< Аa�    XOS�  C�/<   /. a���� POJ�gJ�  C�f�p `�  /. a�����XO-@��/. a�����XO-@��f� n�� ( ( I��-@��/. a����XO .��r
�` �x  NV  /9    a���ƐXO @( I�/ a�    XON^NuNV��-I�� . r��   �-@��J. gH��    l" 爐�� |    ���  )�g(/. . I�/ C��� y    N�PO"n�� @ 	"�N^NuJ. f$ .����    l�" 爐�� |    ���  )�f�/<   /. a�����POJ�gp�-@��`$/. a���žXO @( I�-@��/. a����XO. ��J���lp`    p�� ��� . r��   ��� �� . ���   ��� �� . ��   ����. ���� ���  ��/ �����  ��/ �� ���  ��/ /.��/<  e�a�    ��  N���� ` ��NV  / .  |    "p  	gr (q  g
�  $B� �R��   m�(_N^NuNV  ///(|    B�    `     L�� �  )�gR�     9    ��    m� 9    ��    m/<  e�a�    XO*|    B�    `     M�� �  )�gR�     9    ��    m� 9    ��    m/<  e�a�    XO�� �    @ fnr���    fd 9    r� |   ���  ��t� |   ��  �  ��ኂ���!   �  ��銂���    �  ����� �����#�    J�    gt��    #�  ;�     y    N�$(_*_N^NuNV  #�        #�  ;�    #�        #�  :H    B�    B�    #�  =�    N^NuNV��//*n   |    -p ��g n��p�( $g
p(_*_N^Nu r� �/   -@��B��� .��ሀ���-@��/ a�����XO-@��g  MX�".�� �Ё��� �����`  �    /.��a���XO(@ MX�".�� �Ё����� � �   �!@  MX�".�� �Ё��� � /<   Hl  MX�".�� �Ё���Hh a�    ��  MX�".�� �Ё���B( /<   Hl & MX�".�� �Ё���Hh a�    ��  MX�".�� �Ё���B(  /.��a����XOR���p����n ��p�+@ p ` ��    >A.�&֕5���NqNq      �   2  �  C�  C�  C�  D  D  D  D/  D>  DK  DW  Dg  Dt  D�  D�  D�  D�    D�   D�   D�   E   E   E9   EN   Ee   E�   E�   E�   E�   F   F1   FB  F`  Fq   F�  F�  F�  G  G7   Gb   G�   G�   G�  G�  H	   H=	  HS	  Hj	  H~
   H�   H�  H�  H�   I   I  I2  II  Ic  Ix  I�  I�  I�  I�	  J
  J  J+  J[   J�   J�   J�  J�  K  K"  K8   KM  Kf  K�   K�   K�  L   L  LE  Ln  L�  L�  L�   M,  MY  M�  M�  M�  M�   N  N#  N=  N_   N   N�   N�  N�  N�   O   O.    OO!   On!  O�"   O�$   O�%   O�&   O�&  P
&  P"&  P:'   P](   Pn(  P�)   P�*   P�*  Q	*  Q!+   Q8,   Qi,  Q�,  Q�-   Q�/   Q�0   R0  R+0  RO0  Rx1   R�1  R�2   R�2  R�3   S6   S7   S19   SC:   Sc;   Sv;  S�;  S�;  S�;  T;  T!;  T+;  TG;  Tf;	  Tw;
  T�;  T�;  T�;  T�;  U=   U'>   UH?   Uq?  U�?  U�?  U�@   U�@�  U�A   V!B   V3C   VQD   V_E   VwF   V�G   V�H   V�I   V�J   V�K   WL   W!N   WHP   WfP  WyP  W�Q   W�R   W�S  W�S  W�S   XT   XU   XBW   XZX   X~Y   X�Z   X�Z   X�Z   X�Z   Y[   Y1[   Y?[   YW[   Yn\   Y�\  Y�\  Y�`   Y�a   Y�a  Y�a  Zb   Zc   Z/d   ZZ        No Sense Recovered Error Not Ready Medium Error Hardware Error Illegal Request Unit Attention Data Protect Blank Check Vendor Specific Copy Aborted Aborted Command Equal Volume Overflow Miscompare Reserved No Additional Sense Information Filemark Detected End-Of-Partition/Medium Detected Setmark Detected Beginning-Of-Partition/Medium Detected End-Of-Data Detected I/O Process Terminated Audio Play Operation In Progress Audio Play Operation Paused Audio Play Operation Successfully Completed Audio Play Operation Stopped Due To Error No Current Audio Status To Return No Index/Sector Signal No Seek Complete Peripheral Device Write Fault No Write Current Excessive Write Errors Logical Unit Not Ready Logical Unit Is In Proces Of Becomming Ready Logical Unit Not Ready, Initializing Command Required Logical Unit Not Ready, Manual Intervention Required Logical Unit Not Ready, Format In Progress Logical Unit Does Not Respond To Selection No Reference Position Found Multiple Peripheral Devices Selected Logical Unit Communication Failure Logical Unit Communication Time-Out Logical Unit Communication Parity Error Track Following Error Tracking Servo Failure Focus Servo Failure Spindle Servo Failure Error Log Overflow Write Error Write Error Recovered With Auto-Reallocation Write Error - Auto-Reallocation Failed ID CRC or ECC Error Unrecovered Read Error Read Retries Exhausted Error Too Long To Correct Multiple Read Errors Unrecovered Read Error - Auto-Reallocate Failed L-EC Uncorrectable Error CIRC Unrecovered Error Data Resynchronization Error Incomplete Block Read No Gap Found Miscorrected Error Unrecovered Read Error - Recommend Reassignment Unrecovered Read Error - Recommend Rewrite The Data Address Mark Not Found For ID Field Address Mark Not Found For Data Field Recorded Entity Not Found Record Not Found Filemark Or Setmark Not Found End-Of-Data Not Found Block Sequence Error Random Positioning Error Mechanical Positioning Error Positioning Error Detected By Read Of Medium Data Synchronization Mark Error Recovered Data With No Error Correction Applied Recovered Data With Retries Recovered Data With Positive Head Offset Recovered Data With Negative Head Offset Recovered Data With Retries And/Or CIRC Applied Recovered Data Using Previous Sector ID Recovered Data Without ECC - Data Auto-Reallocated Recovered Data Without ECC - Recommed Reassignment Recovered Data With Error Correction Applied Recovered Data With Error Correction And Retries Applied Recovered Data - Data Auto-Reallocated Recovered Data With CIRC Recovered Data With LEC Recovered Data - Recommed Reassignment Defect List Error Defect List Not Available Defect List Error In Primary List Defect List Error In Grown List Parameter List Length Error Synchronous Data Transfer Error Defect List Not Found Primary Defect List Not Found Grown Defect List Not Found Miscompare During Verify Operation Recovered ID With ECC Correction Invalid Command Operation Code Logical Block Address Out Of Range Invalid Element Address Illegal Function Invalid Field in CDB Logical Unit Not Supported Invalid Field In Parameter List Parameter Not Supported Parameter Value Invalid Threshold Parameters Not Supported Write Protected  Not Ready To Ready Transition (Medium May Have Changed) Import Or Export Element Accessed Power On, Reset, or Bus Device Reset Occurred Parameters Changed Mode Parameters Changed Log Parameters Changed Copy Cannot Execute Since Host Cannot Disconnect Command Sequence Error Too Many Windows Specified Invalid Combination Of Windows Specified Overwrite Error On Update In Place Commands Cleared By Another Initiator Incompatible Medium Installed Cannot Read Medium - Unknown Format Cannot Read Medium - Incompatible Format Cleaning Cartridge Installed Medium Format Corrupted Format Command Failed No Defect Spare Location Available Defect List Update Failure Tape Length Error Ribbon, Ink, or Toner Failure Rounded Parameter Saving Parameters Not Supported Medium Not Present Sequential Positioning Error Tape Position Error At Beginning-Of-Medium Tape Position Error At End-Of-Medium Tape Or Electronic Vertical Forms Unit Not Ready Slew Failure Paper Jam Failed To Sense Top-Of-Form Failed To Sense Bottom-Of-Form Reposition Error Read Past End Of Medium Read Past Beginning Of Medium Position Past End Of Medium Position Past Beginning Of Medium Medium Destination Element Full Medium Source Element Empty Invalid Bits In Identify Message Logical Unit Has Not Self-Configured Yet Target Operating Conditions Have Changed Microcode Has Been Changed Change Operating Definition Inquiry Data Has Changed RAM Failure Diagnostic Failure On Component NN (80-FF) Data Path Failure Power-On or Self-Test Failure Message Error Internal Target Failure Select or Reselect Failure Unsuccessful Soft Reset SCSI Parity Error Initiator Detected Error Message Received Invalid Message Error Command Phase Error Data Phase Error Logical Unit Failed Self-Configuration Overlapped Commands Attempted Write Append Error Write Append Position Error Position Error Related To Timing Erase Failure Cartridge Fault Media Load or Eject Failed Unload Tape Failure Medium Removal Prevented SCSI To Host System Interface Failure System Resource Failure Unable To Recover Table-Of-Contents Generation Does Not Exist Updated Block Read Operator Request or State Change Input Operator Medium Removal Request Operator Selected Write Protect Operator Selected Write Permit Log Exception Threshold Condition Met Log Counter At Maximum Log List Codes Exhausted RPL Status Change Spindles Synchronized Spindles Not Synchronized Lamp Failure Video Acquisition Error Unable To Acquire Video Out Of Focus Scan Head Positioning Error End Of User Area Encountered On This Track Illegal Mode For This Track SCSI: %s
 	(%s)
 major(dev) != 0xff && minor(dev) != 0xffffff ../s200io/scsi.c major(dev) == scsi_blk_major || major(dev) == scsi_raw_major ../s200io/scsi.c (unsigned)m_selcode(dev) < MAX_SCSI_SELCODE ../s200io/scsi.c scsi_card[m_selcode(dev)] != NULL ../s200io/scsi.c scsi_card[m_selcode(dev)]->dev[m_busaddr(dev)] != NULL ../s200io/scsi.c scsi_card[m_selcode(dev)]->dev[m_busaddr(dev)] 		->lun[m_unit(dev)] != NULL ../s200io/scsi.c %s%02x   
	 
 scsi_teac_read
  SCSI: dev = 0x%x: Power On, Reset, or Bus Device Reset Occurred
 SCSI: dev = 0x%x, offset = 0x%x, bcount = 0x%x  b_flags = 0x%x
 	sense key = 0x%x, code = 0x%x, qualifier = 0x%x , info = 0x%x 
 	hexadecimal sense dump:
	 SCSI: deferred error
 SCSI: CDROM: deferred error
 SCSI: unrecoverable deferred error
 	key = 0x%x, code = 0x%x
 SCSI: unrecoverable deferred error un SCSI: %s%s recoverable I/O error  on dev 0x%x at lba 0x%x
 SCSI: scsi_cmd: %d-byte cmd; cmd_mode = 0x%x; clock_ticks = %d: SCSI: disconnect timed out; dev = 0x%x
 SCSI: request timed out; dev = 0x%x; state = 0x%x
 SCSI: select timed out; dev = 0x%x
 FSM: dev = 0x%x, state = 0x%x
 Select (%d): not owner
 scsi: no device at %x
 scsi: select cmd timed out %x
 SCSI mesg in: save_data_ptr
 SCSI mesg in: restore_ptr
 SCSI mesg in: no_op
 SCSI mesg in: disconnect
 SCSI mesg in: Msg Reject
 SCSI: sync negotiation rejected
 SCSI Unknown msg reject (dev: %x)
 SCSI mesg in: cmd complete
 SCSI_SANITY: %s
 MSGcmd_complete SCSI: Bad status from sense
 SCSI: inconsistency in sense
 SCSI: b_error = %d
 SCSI: extended mesg
 SCSI: sync xfr enabled: (io_sync = 0x%x)
 SCSI: unexpected msg: SCSI mesg in: identify %x
 SCSI FSM: Unknown msg_in byte: %x
 SCSI_SANITY: %s
 phase_cmd SCSI_SANITY: %s
 data in / out SCSI data xfr count: %x addr: 0x%x
 SCSI_SANITY: %s
 phase_status SCSI: bad status = 0x%x
 SCSI: Unknown state = 0x%x, phase = 0x%x,  iob->io_sanity = 0x%x
 SCSI: recover: dev = 0x%x, escapecode = %d
 	offset = 0x%x, bcount = 0x%x
 SCSI: scsi_if_abort failed; dev = 0x%x
 unknown state in driver ctl SCSI: dev = 0x%x; inquiry data: SCSI: dev 0x%x has %d %d-byte blocks
 M_IOSYS < M_LAST ../s200io/scsi.c BUCKETINDX(sizeof(*(cp))) <= MAXBUCKET ../s200io/scsi.c M_IOSYS < M_LAST ../s200io/scsi.c BUCKETINDX(sizeof(*(dp))) <= MAXBUCKET ../s200io/scsi.c M_IOSYS < M_LAST ../s200io/scsi.c BUCKETINDX(sizeof(*(up))) <= MAXBUCKET ../s200io/scsi.c  M_IOSYS < M_LAST ../s200io/scsi.c kalloc_aligned((unsigned long)up) ../s200io/scsi.c kup->ku_pagecnt == 0 ../s200io/scsi.c  M_IOSYS < M_LAST ../s200io/scsi.c kalloc_aligned((unsigned long)dp) ../s200io/scsi.c kup->ku_pagecnt == 0 ../s200io/scsi.c  M_IOSYS < M_LAST ../s200io/scsi.c kalloc_aligned((unsigned long)cp) ../s200io/scsi.c kup->ku_pagecnt == 0 ../s200io/scsi.c TEAC     FC-1     HF   07 FC-1     HF   00 !(bp->b_flags & B_DONE) ../s200io/scsi.c MSUS: log2blk %x sc %x unit %x ba %x
 scsi_init: scsi_open not in bdevsw scsi_init: scsi_open not in cdevsw         
  0 _isc_table   �    _cnt   �    _rate   �    _sum   8    _total       _nswap      0 _rootdev       _swapdev       _swapdev_vp    
   _argdev_vp       _nswdev       _mpid       _kmapwnt       _updlock       _rablock       _rasize       _physmembase       _p1pages    
   _highpages    	   _usrstack    
   _user_area       _float_area    
   _processor       _total_lockable_mem       _lockable_mem       _unlockable_mem       _float_present       _dragon_present      0 _bdevsw      0 _cdevsw   (    _linesw   $    _swdevt       _dma32_chan0       _dma32_chan1    	   _dma_here       _free_dma_channels    	   _dmachain   T    _dmatab       _bus_master_count     
   _rupttable   $    _cp_time       0 _dk_devt      0 _dk_busy       0 _dk_time       0 _dk_seek       0 _dk_xfer       0 _dk_wds       0 _dk_mspw       _tk_nin       _tk_nout  ?#   _scsi_max_retries      0 _scsi_bp_lock      0 _scsi_ctl_bp  ?#   _SELECT_TICKS  ? #   _WATCHDOG_TICKS  ?$#   _DISCONNECT_TICKS   � 
  0 _scsi_card      0 _scsi_blk_major      0 _scsi_raw_major  ?(#   _scsi_sense_key  ?h#   _scsi_as    "   _decode_opcode        _msg_printf   �"
   _m_scsi_up       0 _assertions        _assfail  �"   _msg_hex_dmp  "   _scsi_teac_read       0 _SCSI_DEBUG        _ten_byte_cmd  �"   _scsi_decode_sense        _panic  �"	   _scsi_cmd        _scsi_if_transfer  >"   _scsi_discon_timedout        _scsi_if_remove_busfree       0 _fhs_timeout_proc       0 _scsi_if_dequeue        _sw_trigger       0 _flag_timeout  �"   _scsi_req_timedout  	�"   _scsi_select_timedout        _scsi_if_term_arbit  
b"   _scsi_dequeue  
�"	   _scsi_fsm        _C__tst        _C__try        _clear_timeout        _escape        _get_selcode        _C__rec     	   _Ktimeout        _scsi_if_select        _drop_selcode        _scsi_if_clear_reselect     
   _queuedone        _scsi_set_state        _set_smart_poll        _scsi_if_wait_for_reselect       0 _scsi_xfer_cmd       0 _scsi_request_sense       0 _scsi_short_xfer_cmd        ___float        ___fmul        ___dtof        _scsi_if_request_sync_data        _scsi_if_mesg_out        _hidden_mode_exists        _scsi_if_status        _scsi_if_mesg_in       0 _u        _scsi_if_abort  F"	   _scsi_nop  Z"   _scsi_driver_ctl        _enqueue       0 _scsi_start_stop       0 _scsi_move_medium       0 _scsi_init_element_status       0 _scsi_read_element_status       0 _scsi_reserve       0 _scsi_release  �"   _scsi_control       0 _scsi_format_unit        _geteblk        _sleep       0 _scsi_mode_select        _bcopy        _biowait       0 _scsi_inquiry       0 _scsi_read_capacity        _brelse        _wakeup     	   _geterror  |"   _scsi_lun_open       0 _bucket        _CRIT       0 _mpproc_info     	  0 _kmemlock        _UNCRIT        _kmalloc     
  0 _kmemstats        _bzero  #�"   _scsi_lun_close     
   _page_info        _kalloc_aligned        _kfree  C�#   _flush_on_all_closes  (�"   _scsi_close     
   _sds_close  -"   _scsi_free_dk_index        _dma_unactive       0 _scsi_allow_media  )�"
   _scsi_open     	   _sds_open  ,~"   _scsi_assign_dk_index        _dma_active        _strncmp       0 _scsi_test_unit  0l"   _scsi_init_capacity       0 _scsi_prevent_media  -<"   _scsi_teac_setup       0 _scsi_mode_sense_cmd  .�"   _scsi_teac_init_capacity  16"   _scsi_ioctl     
   _sds_ioctl        _suser  7V"   _scsi_strategy        _sds_strategy        _biodone        _bpcheck       0 _led_activity_bits  8�"   _scsi_write     
   _sds_write       0 _minphys        _physio  9,"
   _scsi_read     	   _sds_read  9x"
   _scsi_size     	   _sds_size        _snooze  : "
   _scsi_dump       0 _dumpdev        _scsi_if_dump      0 _scsi_saved_msus_for_boot      0 _scsi_saved_dev_init  :H"   _scsi_msus_for_boot       0 _nblkdev       0 _nchrdev  ;�"   _scsi_reset  ;�"
   _scsi_init       0 _msus       0 _striped_boot       0 _scsi_reset_callback  =N"
   _scsi_link     	  0 _dev_init       0 _msus_for_boot  =�"   _scsi_config_identify       0 _scsi_config_ident        _strncpy        _strncat        (     . >   P     n     �     �     � >   � @   �          A   @  $ 9  8 :  F    L    R A  \ @  ~    �    � A  � @  � 8  �    �    � A  � @  � 8      
     A   @  . 8  \    b    h A  ~ 8  �    �    �    � >  �      >  ( D  6    < >  � E  �    F    L >  j    p >  �    � >  �    � >  �    � >  �    � >  �    � >  "    ( >  D    J >  Z    ` >  ~    � >  �    � G  �     �     �     �     �     �     �     �     �     �     �     �     �     H     R    p    z    � >  �    � >  � D  �    � >  � D  , I  P    V >  ` K  � L  � M  � N  � O  	    	 >  	J L  	l M  	v N  	� O  	�    	� >  	� R  	� L  
  M  
* N  
V O  
~ M  
� N  
� U  
� V  
� D       >  * W  B X  �     � Y  � X  � Z  �    �     � [  � \  � W   X  $ D  <    B >  Z ]  n D  �    � >  � ^  � _  �    � >  � X  � ^  � X  $ `  4     : a  J D  Z    ` >  r D  �    � >  � D  �    � >  � D  �    � >  �     � b       
 [   D  (    . >  ^ D  n    t >  � D  �    � >  � *  � c  � .  � D  �    � >      "    ( >  6 X  f    l >  z X  � d  � e  �     ]  "     ( [  ` d  j    p >  �    � ]  � ]   D      $ >  . _  r D  �    � >  �     �     � f  � g  � h  � /   D  $    * >  :    @ >  n D  �    � >  �    � >  � X  � *  � c  � -   ,  " e  � i  �          [   j  ( W  @ X  ^ X  ~    �    � >  � X  �    �     � [  �    �    � >   X   D  (    . >  <    D     J [  n k  z c  � I  � e  �    �    � >   X  &    .     4 [  @ l  \ W  t X  � D  �    � >  � X  �    � >  �    � >   X  �    �     � [  � m  � W  � X  "     (     ,     0     4     8     <     @     D     H     V W  b n  n    t >  �    � >  � *  � ^  � o  �    � >  � ]  � n  0 _  P _  �    �     �     �     �     �     �     �                 r  &     @ s  J t  f u  � v  � w  � x  �    � G  � z  � {  � 3   3   3   |   3  " 4  0 {  8 4  > 4  �    � }  � ~  � r      }  8 ~  B �  X D  f    l >  � �  � ~  � ~  � D  
     >  2 z  > �  J 3  X 3  ^ �  f 3  n �  � 8  � 8  � �  � �  � �  � �   �   �  * �  @ �  R �  � �  � �  � �  � 8  � �  � �    8   6 8   @ |   T 8   � �   � �   � �   � �   � �   � �   � �   � �  ! �  !j �  !v �  !� �  !� �  !� �  !� |  ", �  "4 �  "< �  "\ �  "l �  "x �  "� �  "� �  "� �  # �  # �  #8 �  #R �  #b �  #� |  $ 8  $v �  $� @  $� �  $�    $�    $� A  $� �  $� �  $� �  $� @  %    %    %  A  %* �  %2 �  %R �  %� �  %� �  %� �  %� �  %� @  %� �  &    &    & A  &0 �  &P �  &\ �  &d @  &|    &�    &� A  &� �  &� �  &� �  &� �  ' �  ' �  '> 8  'J �  'V @  'b �  't    'z    '� A  '� �  '� �  '� �  '� @  '�    '�    '� A  '� �  ( �  (" �  (^ �  (j �  (� �  (� �  (�    (�     )6    )@ �  )T :  )� �  )�     )� �  *    *� :  *� �  *� �  *�     +0    +: �  +N    +X �  +l    +v �  +� 9  +�     +�     +�     +�     +�     +�     +�     +�     +�     , �  ,"     ,d �  ,j     ,� )  ,� *  ,� +  ,� -  ,� ,  ,� /  ,�     ,� 9  -  )  -* )  -v �  -|     -� �  -� ~  .p }  .v     /     /$     /t     /z     /�     /�     04     0:     0� �  0�     1 �  1     1` �  1� ~  2� �  2� �  3� ~  3� ~  3� �  4 �  4H     4P     4T     4X     4\     4`     4d     4h     4l     4p     4t     4x     4|     4�     4�     4�     4�     4�     5Z z  5`     5� �  5�     6 �  6     6P ~  7j @  7�    7�    7� A  7� �  7�    7�    7�     8 :  88     8f �  8� �  8� e  8� c  8� �  8� �  8� r  8� �  9 �  9     9" �  9F �  9V �  9h     9n �  9� �  9� �  9�    9�    :& �  :> �  :j �  :z   :�     :� �  :� �  :�   :�     ;�    ;� >  ;� 8  <   < 9  <      <( 9  <. 9  <4 �  << 9  <B �  <J    <P G  <X   <^ :  <p     <x :  <~ :  <� �  <� :  <� �  <�    <� G  <� �  <�   <� 9  <� �  <� �  <� �  = �  =   =$ �  =.   =4     =8 �  => �  =T �  =X �  =^     =b �  =h �  =l �  =r     =v �  =| 3  =� 4  =�     =� �  =�    >� �  >� �                             $     (     ,     0     4     8     <     @     D     H     L     R     X     ^     d     j     p     v     |     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �     �                             $    *    0    6    <    B    H    N    T    Z    `    f    l    r    x    ~    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �                             &    ,    2    8    >    D    J    P    V    \    b    h    n    t    z    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �        
                "    (    .    4    :    @    F    L    R    X    ^    d    j    p    v    |    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �    �                             $    *    0    6    <    B    H    N    T    Z    `    f    l    r    x    ~    �    �    �    �    �    �    �    �    �    �  